/* Test bench for vga_620x480.v
 saved in vga_620x480_tb.v */

`timescale 1ns / 1ps

`include "vga_620x480.v"



module vga_tb;

   reg         clk;
   reg  [15:0] pixel;
   wire        v_sync;
   wire        h_sync;
   wire [3:0]  Red;
   wire [3:0]  Green;
   wire [3:0]  Blue;
   wire [31:0] pixel_ADDR;
   
   // wrapper
   vga UUT(
	   clk,
	   pixel,
	   v_sync,
	   h_sync,
	   Red,
	   Green,
	   Blue,
	   pixel_ADDR
	   );

   // Generate Clock
   initial begin
      clk = 1;
      forever #5 clk = ~clk;
   end

   // Pass pixel address to value for simulation
   initial begin
      forever
	 #10 pixel <= pixel_ADDR[19:4];
   end
   
   
   // Generate Dumpfile and define runtime
   initial begin
      $dumpfile("vga.vcd");
      $dumpvars(0, vga_tb);

      #1000000 $finish;
      
      //#100000000 $finish;
      
   end
   
   

endmodule // vga_tb
